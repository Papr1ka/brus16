

module example_rom_gpu (
    input wire clk,
    input wire[15:0] addr_a, // read only addr
    output reg[15:0] dout_a, // a data
    input wire we_b, // write enable on b
    input wire[15:0] addr_b, // write only addr
    input wire[15:0] din_b // write only data
);

// test rectangles
initial begin
    // rectangles
    ram[0] = 16'b0000000000000001;
    ram[1] = 16'b0000000000000000;
    ram[2] = 16'b0000000000000000;
    ram[3] = 16'b0000000100000000;
    ram[4] = 16'b0000000100000000;
    ram[5] = 16'b0011100100000000;
    ram[6] = 16'b0000000000000001;
    ram[7] = 16'b0000000000000000;
    ram[8] = 16'b0000000000000000;
    ram[9] = 16'b0000000011111100;
    ram[10] = 16'b0000000100000000;
    ram[11] = 16'b0000110011001110;
    ram[12] = 16'b0000000000000001;
    ram[13] = 16'b0000000000000000;
    ram[14] = 16'b0000000000000000;
    ram[15] = 16'b0000000011111000;
    ram[16] = 16'b0000000100000000;
    ram[17] = 16'b1000110011010000;
    ram[18] = 16'b0000000000000001;
    ram[19] = 16'b0000000000000000;
    ram[20] = 16'b0000000000000000;
    ram[21] = 16'b0000000011110100;
    ram[22] = 16'b0000000100000000;
    ram[23] = 16'b0111110101100010;
    ram[24] = 16'b0000000000000001;
    ram[25] = 16'b0000000000000000;
    ram[26] = 16'b0000000000000000;
    ram[27] = 16'b0000000011110000;
    ram[28] = 16'b0000000100000000;
    ram[29] = 16'b0111001001001000;
    ram[30] = 16'b0000000000000001;
    ram[31] = 16'b0000000000000000;
    ram[32] = 16'b0000000000000000;
    ram[33] = 16'b0000000011101100;
    ram[34] = 16'b0000000100000000;
    ram[35] = 16'b0100011101110001;
    ram[36] = 16'b0000000000000001;
    ram[37] = 16'b0000000000000000;
    ram[38] = 16'b0000000000000000;
    ram[39] = 16'b0000000011101000;
    ram[40] = 16'b0000000100000000;
    ram[41] = 16'b0011010001111010;
    ram[42] = 16'b0000000000000001;
    ram[43] = 16'b0000000000000000;
    ram[44] = 16'b0000000000000000;
    ram[45] = 16'b0000000011100100;
    ram[46] = 16'b0000000100000000;
    ram[47] = 16'b0010110010000011;
    ram[48] = 16'b0000000000000001;
    ram[49] = 16'b0000000000000000;
    ram[50] = 16'b0000000000000000;
    ram[51] = 16'b0000000011100000;
    ram[52] = 16'b0000000100000000;
    ram[53] = 16'b1101100000000110;
    ram[54] = 16'b0000000000000001;
    ram[55] = 16'b0000000000000000;
    ram[56] = 16'b0000000000000000;
    ram[57] = 16'b0000000011011100;
    ram[58] = 16'b0000000100000000;
    ram[59] = 16'b0001000001000101;
    ram[60] = 16'b0000000000000001;
    ram[61] = 16'b0000000000000000;
    ram[62] = 16'b0000000000000000;
    ram[63] = 16'b0000000011011000;
    ram[64] = 16'b0000000100000000;
    ram[65] = 16'b0000111101000001;
    ram[66] = 16'b0000000000000001;
    ram[67] = 16'b0000000000000000;
    ram[68] = 16'b0000000000000000;
    ram[69] = 16'b0000000011010100;
    ram[70] = 16'b0000000100000000;
    ram[71] = 16'b0010111111111000;
    ram[72] = 16'b0000000000000001;
    ram[73] = 16'b0000000000000000;
    ram[74] = 16'b0000000000000000;
    ram[75] = 16'b0000000011010000;
    ram[76] = 16'b0000000100000000;
    ram[77] = 16'b0110111111110001;
    ram[78] = 16'b0000000000000001;
    ram[79] = 16'b0000000000000000;
    ram[80] = 16'b0000000000000000;
    ram[81] = 16'b0000000011001100;
    ram[82] = 16'b0000000100000000;
    ram[83] = 16'b0111011100011111;
    ram[84] = 16'b0000000000000001;
    ram[85] = 16'b0000000000000000;
    ram[86] = 16'b0000000000000000;
    ram[87] = 16'b0000000011001000;
    ram[88] = 16'b0000000100000000;
    ram[89] = 16'b0000110110010110;
    ram[90] = 16'b0000000000000001;
    ram[91] = 16'b0000000000000000;
    ram[92] = 16'b0000000000000000;
    ram[93] = 16'b0000000011000100;
    ram[94] = 16'b0000000100000000;
    ram[95] = 16'b0110010111001110;
    ram[96] = 16'b0000000000000001;
    ram[97] = 16'b0000000000000000;
    ram[98] = 16'b0000000000000000;
    ram[99] = 16'b0000000011000000;
    ram[100] = 16'b0000000100000000;
    ram[101] = 16'b1101011011001011;
    ram[102] = 16'b0000000000000001;
    ram[103] = 16'b0000000000000000;
    ram[104] = 16'b0000000000000000;
    ram[105] = 16'b0000000010111100;
    ram[106] = 16'b0000000100000000;
    ram[107] = 16'b0111000011011101;
    ram[108] = 16'b0000000000000001;
    ram[109] = 16'b0000000000000000;
    ram[110] = 16'b0000000000000000;
    ram[111] = 16'b0000000010111000;
    ram[112] = 16'b0000000100000000;
    ram[113] = 16'b1110010111111110;
    ram[114] = 16'b0000000000000001;
    ram[115] = 16'b0000000000000000;
    ram[116] = 16'b0000000000000000;
    ram[117] = 16'b0000000010110100;
    ram[118] = 16'b0000000100000000;
    ram[119] = 16'b1000111001101111;
    ram[120] = 16'b0000000000000001;
    ram[121] = 16'b0000000000000000;
    ram[122] = 16'b0000000000000000;
    ram[123] = 16'b0000000010110000;
    ram[124] = 16'b0000000100000000;
    ram[125] = 16'b0000001101010011;
    ram[126] = 16'b0000000000000001;
    ram[127] = 16'b0000000000000000;
    ram[128] = 16'b0000000000000000;
    ram[129] = 16'b0000000010101100;
    ram[130] = 16'b0000000100000000;
    ram[131] = 16'b0101000110111110;
    ram[132] = 16'b0000000000000001;
    ram[133] = 16'b0000000000000000;
    ram[134] = 16'b0000000000000000;
    ram[135] = 16'b0000000010101000;
    ram[136] = 16'b0000000100000000;
    ram[137] = 16'b1101100001100000;
    ram[138] = 16'b0000000000000001;
    ram[139] = 16'b0000000000000000;
    ram[140] = 16'b0000000000000000;
    ram[141] = 16'b0000000010100100;
    ram[142] = 16'b0000000100000000;
    ram[143] = 16'b1010111000110101;
    ram[144] = 16'b0000000000000001;
    ram[145] = 16'b0000000000000000;
    ram[146] = 16'b0000000000000000;
    ram[147] = 16'b0000000010100000;
    ram[148] = 16'b0000000100000000;
    ram[149] = 16'b1000111001000101;
    ram[150] = 16'b0000000000000001;
    ram[151] = 16'b0000000000000000;
    ram[152] = 16'b0000000000000000;
    ram[153] = 16'b0000000010011100;
    ram[154] = 16'b0000000100000000;
    ram[155] = 16'b0100111110011011;
    ram[156] = 16'b0000000000000001;
    ram[157] = 16'b0000000000000000;
    ram[158] = 16'b0000000000000000;
    ram[159] = 16'b0000000010011000;
    ram[160] = 16'b0000000100000000;
    ram[161] = 16'b0110111000111101;
    ram[162] = 16'b0000000000000001;
    ram[163] = 16'b0000000000000000;
    ram[164] = 16'b0000000000000000;
    ram[165] = 16'b0000000010010100;
    ram[166] = 16'b0000000100000000;
    ram[167] = 16'b1010110001010110;
    ram[168] = 16'b0000000000000001;
    ram[169] = 16'b0000000000000000;
    ram[170] = 16'b0000000000000000;
    ram[171] = 16'b0000000010010000;
    ram[172] = 16'b0000000100000000;
    ram[173] = 16'b0011010001010100;
    ram[174] = 16'b0000000000000001;
    ram[175] = 16'b0000000000000000;
    ram[176] = 16'b0000000000000000;
    ram[177] = 16'b0000000010001100;
    ram[178] = 16'b0000000100000000;
    ram[179] = 16'b0010111101111100;
    ram[180] = 16'b0000000000000001;
    ram[181] = 16'b0000000000000000;
    ram[182] = 16'b0000000000000000;
    ram[183] = 16'b0000000010001000;
    ram[184] = 16'b0000000100000000;
    ram[185] = 16'b1100001010000101;
    ram[186] = 16'b0000000000000001;
    ram[187] = 16'b0000000000000000;
    ram[188] = 16'b0000000000000000;
    ram[189] = 16'b0000000010000100;
    ram[190] = 16'b0000000100000000;
    ram[191] = 16'b0011000110000100;
    ram[192] = 16'b0000000000000001;
    ram[193] = 16'b0000000000000000;
    ram[194] = 16'b0000000000000000;
    ram[195] = 16'b0000000010000000;
    ram[196] = 16'b0000000100000000;
    ram[197] = 16'b1011011111001100;
    ram[198] = 16'b0000000000000001;
    ram[199] = 16'b0000000000000000;
    ram[200] = 16'b0000000000000000;
    ram[201] = 16'b0000000001111100;
    ram[202] = 16'b0000000100000000;
    ram[203] = 16'b1011000000011010;
    ram[204] = 16'b0000000000000001;
    ram[205] = 16'b0000000000000000;
    ram[206] = 16'b0000000000000000;
    ram[207] = 16'b0000000001111000;
    ram[208] = 16'b0000000100000000;
    ram[209] = 16'b1000011101101111;
    ram[210] = 16'b0000000000000001;
    ram[211] = 16'b0000000000000000;
    ram[212] = 16'b0000000000000000;
    ram[213] = 16'b0000000001110100;
    ram[214] = 16'b0000000100000000;
    ram[215] = 16'b0001011000111111;
    ram[216] = 16'b0000000000000001;
    ram[217] = 16'b0000000000000000;
    ram[218] = 16'b0000000000000000;
    ram[219] = 16'b0000000001110000;
    ram[220] = 16'b0000000100000000;
    ram[221] = 16'b1110101100111001;
    ram[222] = 16'b0000000000000001;
    ram[223] = 16'b0000000000000000;
    ram[224] = 16'b0000000000000000;
    ram[225] = 16'b0000000001101100;
    ram[226] = 16'b0000000100000000;
    ram[227] = 16'b0011111111101001;
    ram[228] = 16'b0000000000000001;
    ram[229] = 16'b0000000000000000;
    ram[230] = 16'b0000000000000000;
    ram[231] = 16'b0000000001101000;
    ram[232] = 16'b0000000100000000;
    ram[233] = 16'b1100000111001111;
    ram[234] = 16'b0000000000000001;
    ram[235] = 16'b0000000000000000;
    ram[236] = 16'b0000000000000000;
    ram[237] = 16'b0000000001100100;
    ram[238] = 16'b0000000100000000;
    ram[239] = 16'b0010100001011000;
    ram[240] = 16'b0000000000000001;
    ram[241] = 16'b0000000000000000;
    ram[242] = 16'b0000000000000000;
    ram[243] = 16'b0000000001100000;
    ram[244] = 16'b0000000100000000;
    ram[245] = 16'b1001011000011011;
    ram[246] = 16'b0000000000000001;
    ram[247] = 16'b0000000000000000;
    ram[248] = 16'b0000000000000000;
    ram[249] = 16'b0000000001011100;
    ram[250] = 16'b0000000100000000;
    ram[251] = 16'b1011100100101000;
    ram[252] = 16'b0000000000000001;
    ram[253] = 16'b0000000000000000;
    ram[254] = 16'b0000000000000000;
    ram[255] = 16'b0000000001011000;
    ram[256] = 16'b0000000100000000;
    ram[257] = 16'b0110001001110011;
    ram[258] = 16'b0000000000000001;
    ram[259] = 16'b0000000000000000;
    ram[260] = 16'b0000000000000000;
    ram[261] = 16'b0000000001010100;
    ram[262] = 16'b0000000100000000;
    ram[263] = 16'b0010001110011100;
    ram[264] = 16'b0000000000000001;
    ram[265] = 16'b0000000000000000;
    ram[266] = 16'b0000000000000000;
    ram[267] = 16'b0000000001010000;
    ram[268] = 16'b0000000100000000;
    ram[269] = 16'b0001011101110110;
    ram[270] = 16'b0000000000000001;
    ram[271] = 16'b0000000000000000;
    ram[272] = 16'b0000000000000000;
    ram[273] = 16'b0000000001001100;
    ram[274] = 16'b0000000100000000;
    ram[275] = 16'b0111010010101111;
    ram[276] = 16'b0000000000000001;
    ram[277] = 16'b0000000000000000;
    ram[278] = 16'b0000000000000000;
    ram[279] = 16'b0000000001001000;
    ram[280] = 16'b0000000100000000;
    ram[281] = 16'b1001010000101010;
    ram[282] = 16'b0000000000000001;
    ram[283] = 16'b0000000000000000;
    ram[284] = 16'b0000000000000000;
    ram[285] = 16'b0000000001000100;
    ram[286] = 16'b0000000100000000;
    ram[287] = 16'b0010100011011010;
    ram[288] = 16'b0000000000000001;
    ram[289] = 16'b0000000000000000;
    ram[290] = 16'b0000000000000000;
    ram[291] = 16'b0000000001000000;
    ram[292] = 16'b0000000100000000;
    ram[293] = 16'b0111011100110000;
    ram[294] = 16'b0000000000000001;
    ram[295] = 16'b0000000000000000;
    ram[296] = 16'b0000000000000000;
    ram[297] = 16'b0000000000111100;
    ram[298] = 16'b0000000100000000;
    ram[299] = 16'b0011001110110110;
    ram[300] = 16'b0000000000000001;
    ram[301] = 16'b0000000000000000;
    ram[302] = 16'b0000000000000000;
    ram[303] = 16'b0000000000111000;
    ram[304] = 16'b0000000100000000;
    ram[305] = 16'b1100001010011111;
    ram[306] = 16'b0000000000000001;
    ram[307] = 16'b0000000000000000;
    ram[308] = 16'b0000000000000000;
    ram[309] = 16'b0000000000110100;
    ram[310] = 16'b0000000100000000;
    ram[311] = 16'b1000111001010010;
    ram[312] = 16'b0000000000000001;
    ram[313] = 16'b0000000000000000;
    ram[314] = 16'b0000000000000000;
    ram[315] = 16'b0000000000110000;
    ram[316] = 16'b0000000100000000;
    ram[317] = 16'b1110100000100101;
    ram[318] = 16'b0000000000000001;
    ram[319] = 16'b0000000000000000;
    ram[320] = 16'b0000000000000000;
    ram[321] = 16'b0000000000101100;
    ram[322] = 16'b0000000100000000;
    ram[323] = 16'b1011101011001011;
    ram[324] = 16'b0000000000000001;
    ram[325] = 16'b0000000000000000;
    ram[326] = 16'b0000000000000000;
    ram[327] = 16'b0000000000101000;
    ram[328] = 16'b0000000100000000;
    ram[329] = 16'b0101001101000111;
    ram[330] = 16'b0000000000000001;
    ram[331] = 16'b0000000000000000;
    ram[332] = 16'b0000000000000000;
    ram[333] = 16'b0000000000100100;
    ram[334] = 16'b0000000100000000;
    ram[335] = 16'b1011110110001000;
    ram[336] = 16'b0000000000000001;
    ram[337] = 16'b0000000000000000;
    ram[338] = 16'b0000000000000000;
    ram[339] = 16'b0000000000100000;
    ram[340] = 16'b0000000100000000;
    ram[341] = 16'b1011010111100110;
    ram[342] = 16'b0000000000000001;
    ram[343] = 16'b0000000000000000;
    ram[344] = 16'b0000000000000000;
    ram[345] = 16'b0000000000011100;
    ram[346] = 16'b0000000100000000;
    ram[347] = 16'b0110101101000100;
    ram[348] = 16'b0000000000000001;
    ram[349] = 16'b0000000000000000;
    ram[350] = 16'b0000000000000000;
    ram[351] = 16'b0000000000011000;
    ram[352] = 16'b0000000100000000;
    ram[353] = 16'b1000100010110001;
    ram[354] = 16'b0000000000000001;
    ram[355] = 16'b0000000000000000;
    ram[356] = 16'b0000000000000000;
    ram[357] = 16'b0000000000010100;
    ram[358] = 16'b0000000100000000;
    ram[359] = 16'b0010010010001110;
    ram[360] = 16'b0000000000000001;
    ram[361] = 16'b0000000000000000;
    ram[362] = 16'b0000000000000000;
    ram[363] = 16'b0000000000010000;
    ram[364] = 16'b0000000100000000;
    ram[365] = 16'b0101011110011111;
    ram[366] = 16'b0000000000000001;
    ram[367] = 16'b0000000000000000;
    ram[368] = 16'b0000000000000000;
    ram[369] = 16'b0000000000001100;
    ram[370] = 16'b0000000100000000;
    ram[371] = 16'b0111110101010111;
    ram[372] = 16'b0000000000000001;
    ram[373] = 16'b0000000000000000;
    ram[374] = 16'b0000000000000000;
    ram[375] = 16'b0000000000001000;
    ram[376] = 16'b0000000100000000;
    ram[377] = 16'b0101001110101001;
    ram[378] = 16'b0000000000000001;
    ram[379] = 16'b0000000000000000;
    ram[380] = 16'b0000000000000000;
    ram[381] = 16'b0000000000000100;
    ram[382] = 16'b0000000100000000;
    ram[383] = 16'b1110110010101101;
end

reg [15:0] ram [1023:0];

always @(posedge clk) begin
    dout_a <= ram[addr_a[9:0]];
    if (we_b) begin
        ram[addr_b[9:0]] <= din_b;
    end
end

endmodule
