/*
    1*READ 1*WRITE sync memory
    intended to be implemented as block ram
    sync read, sync write
*/
module bsram
#(
    parameter WIDTH = 13,
    parameter SIZE = 8192,
    parameter PROGRAM = 1
)
(
    input wire clk,

    // read
    input wire [WIDTH-1:0] mem_dout_addr,
    output reg [15:0] mem_dout,
    
    // write
    input wire we,
    input wire [WIDTH-1:0] mem_din_addr,
    input wire [15:0] mem_din
);

reg [15:0] data [SIZE-1:0];

always @(posedge clk) begin
    if (we) begin
        data[mem_din_addr] <= mem_din;
    end
    mem_dout <= data[mem_dout_addr];
end

initial begin
    for (integer i = 0; i < SIZE; i = i + 1) begin
        data[i] = 16'b0;
    end
    if (PROGRAM) begin
        // game program
        data[0] = 65140;
        data[1] = 19456;
        data[2] = 49161;
        data[3] = 23041;
        data[4] = 40968;
        data[5] = 49166;
        data[6] = 25600;
        data[7] = 32771;
        data[8] = 22016;
        data[9] = 23286;
        data[10] = 65152;
        data[11] = 57344;
        data[12] = 49662;
        data[13] = 22016;
        data[14] = 49171;
        data[15] = 49235;
        data[16] = 49428;
        data[17] = 49293;
        data[18] = 22016;
        data[19] = 65142;
        data[20] = 16384;
        data[21] = 23552;
        data[22] = 40990;
        data[23] = 57613;
        data[24] = 16384;
        data[25] = 23552;
        data[26] = 522;
        data[27] = 57613;
        data[28] = 17408;
        data[29] = 32798;
        data[30] = 65143;
        data[31] = 16384;
        data[32] = 23552;
        data[33] = 41004;
        data[34] = 57613;
        data[35] = 16384;
        data[36] = 23552;
        data[37] = 1556;
        data[38] = 57613;
        data[39] = 17408;
        data[40] = 23040;
        data[41] = 57612;
        data[42] = 17408;
        data[43] = 32812;
        data[44] = 65140;
        data[45] = 16384;
        data[46] = 23552;
        data[47] = 41018;
        data[48] = 57613;
        data[49] = 16384;
        data[50] = 23552;
        data[51] = 14948;
        data[52] = 41017;
        data[53] = 23522;
        data[54] = 57612;
        data[55] = 17408;
        data[56] = 32825;
        data[57] = 32826;
        data[58] = 65141;
        data[59] = 16384;
        data[60] = 23552;
        data[61] = 41032;
        data[62] = 57613;
        data[63] = 16384;
        data[64] = 23552;
        data[65] = 14948;
        data[66] = 41031;
        data[67] = 23070;
        data[68] = 57612;
        data[69] = 17408;
        data[70] = 32839;
        data[71] = 32840;
        data[72] = 57613;
        data[73] = 16384;
        data[74] = 23552;
        data[75] = 1539;
        data[76] = 23040;
        data[77] = 49632;
        data[78] = 59344;
        data[79] = 49647;
        data[80] = 57613;
        data[81] = 17408;
        data[82] = 22016;
        data[83] = 18946;
        data[84] = 23041;
        data[85] = 59344;
        data[86] = 57613;
        data[87] = 16384;
        data[88] = 23552;
        data[89] = 1024;
        data[90] = 7689;
        data[91] = 0;
        data[92] = 17920;
        data[93] = 57612;
        data[94] = 16384;
        data[95] = 23552;
        data[96] = 13824;
        data[97] = 41069;
        data[98] = 57612;
        data[99] = 16384;
        data[100] = 23552;
        data[101] = 16896;
        data[102] = 23552;
        data[103] = 1024;
        data[104] = 23040;
        data[105] = 49632;
        data[106] = 57612;
        data[107] = 17408;
        data[108] = 32893;
        data[109] = 57612;
        data[110] = 16384;
        data[111] = 23552;
        data[112] = 11776;
        data[113] = 41085;
        data[114] = 57612;
        data[115] = 16384;
        data[116] = 23552;
        data[117] = 16896;
        data[118] = 23552;
        data[119] = 0;
        data[120] = 23040;
        data[121] = 49647;
        data[122] = 57612;
        data[123] = 17408;
        data[124] = 32893;
        data[125] = 65279;
        data[126] = 16384;
        data[127] = 23552;
        data[128] = 17921;
        data[129] = 16897;
        data[130] = 23552;
        data[131] = 57612;
        data[132] = 16384;
        data[133] = 23552;
        data[134] = 516;
        data[135] = 23043;
        data[136] = 8192;
        data[137] = 0;
        data[138] = 65279;
        data[139] = 17408;
        data[140] = 22018;
        data[141] = 18945;
        data[142] = 65314;
        data[143] = 17920;
        data[144] = 16896;
        data[145] = 23552;
        data[146] = 514;
        data[147] = 16384;
        data[148] = 23552;
        data[149] = 58324;
        data[150] = 14336;
        data[151] = 16896;
        data[152] = 23552;
        data[153] = 514;
        data[154] = 16384;
        data[155] = 23552;
        data[156] = 57844;
        data[157] = 3071;
        data[158] = 12288;
        data[159] = 4096;
        data[160] = 41150;
        data[161] = 49695;
        data[162] = 58344;
        data[163] = 15360;
        data[164] = 41149;
        data[165] = 57594;
        data[166] = 49695;
        data[167] = 3587;
        data[168] = 0;
        data[169] = 16384;
        data[170] = 23552;
        data[171] = 16896;
        data[172] = 23552;
        data[173] = 513;
        data[174] = 17408;
        data[175] = 23472;
        data[176] = 16896;
        data[177] = 23552;
        data[178] = 514;
        data[179] = 17408;
        data[180] = 57598;
        data[181] = 49695;
        data[182] = 3587;
        data[183] = 0;
        data[184] = 16384;
        data[185] = 23552;
        data[186] = 57614;
        data[187] = 17408;
        data[188] = 32957;
        data[189] = 32977;
        data[190] = 16896;
        data[191] = 23552;
        data[192] = 514;
        data[193] = 16384;
        data[194] = 23552;
        data[195] = 57614;
        data[196] = 16384;
        data[197] = 23552;
        data[198] = 3071;
        data[199] = 57613;
        data[200] = 16384;
        data[201] = 23552;
        data[202] = 7687;
        data[203] = 0;
        data[204] = 0;
        data[205] = 16896;
        data[206] = 23552;
        data[207] = 514;
        data[208] = 17408;
        data[209] = 65350;
        data[210] = 17920;
        data[211] = 16896;
        data[212] = 23552;
        data[213] = 514;
        data[214] = 16384;
        data[215] = 23552;
        data[216] = 57824;
        data[217] = 14336;
        data[218] = 16896;
        data[219] = 23552;
        data[220] = 514;
        data[221] = 16384;
        data[222] = 23552;
        data[223] = 57844;
        data[224] = 3071;
        data[225] = 12288;
        data[226] = 4096;
        data[227] = 41217;
        data[228] = 49695;
        data[229] = 58344;
        data[230] = 15360;
        data[231] = 41216;
        data[232] = 57602;
        data[233] = 49695;
        data[234] = 3587;
        data[235] = 0;
        data[236] = 16384;
        data[237] = 23552;
        data[238] = 16896;
        data[239] = 23552;
        data[240] = 513;
        data[241] = 17408;
        data[242] = 23352;
        data[243] = 16896;
        data[244] = 23552;
        data[245] = 514;
        data[246] = 17408;
        data[247] = 57606;
        data[248] = 49695;
        data[249] = 3587;
        data[250] = 0;
        data[251] = 16384;
        data[252] = 23552;
        data[253] = 57615;
        data[254] = 17408;
        data[255] = 33024;
        data[256] = 33043;
        data[257] = 16896;
        data[258] = 23552;
        data[259] = 514;
        data[260] = 16384;
        data[261] = 23552;
        data[262] = 57615;
        data[263] = 16384;
        data[264] = 23552;
        data[265] = 57613;
        data[266] = 16384;
        data[267] = 23552;
        data[268] = 7687;
        data[269] = 0;
        data[270] = 0;
        data[271] = 16896;
        data[272] = 23552;
        data[273] = 514;
        data[274] = 17408;
        data[275] = 22017;
        data[276] = 18945;
        data[277] = 57613;
        data[278] = 16384;
        data[279] = 23552;
        data[280] = 7687;
        data[281] = 17920;
        data[282] = 16896;
        data[283] = 23552;
        data[284] = 49574;
        data[285] = 16896;
        data[286] = 23552;
        data[287] = 49449;
        data[288] = 16896;
        data[289] = 23552;
        data[290] = 65230;
        data[291] = 49524;
        data[292] = 16896;
        data[293] = 23552;
        data[294] = 65254;
        data[295] = 49524;
        data[296] = 22017;
        data[297] = 18947;
        data[298] = 17920;
        data[299] = 65200;
        data[300] = 17921;
        data[301] = 65176;
        data[302] = 17922;
        data[303] = 16897;
        data[304] = 23552;
        data[305] = 514;
        data[306] = 16384;
        data[307] = 23552;
        data[308] = 57824;
        data[309] = 14336;
        data[310] = 49695;
        data[311] = 58344;
        data[312] = 15360;
        data[313] = 3072;
        data[314] = 41294;
        data[315] = 16898;
        data[316] = 23552;
        data[317] = 514;
        data[318] = 16384;
        data[319] = 23552;
        data[320] = 11776;
        data[321] = 41293;
        data[322] = 16898;
        data[323] = 23552;
        data[324] = 514;
        data[325] = 16384;
        data[326] = 23552;
        data[327] = 1609;
        data[328] = 16897;
        data[329] = 23552;
        data[330] = 514;
        data[331] = 17408;
        data[332] = 33101;
        data[333] = 33102;
        data[334] = 16897;
        data[335] = 23552;
        data[336] = 514;
        data[337] = 16384;
        data[338] = 23552;
        data[339] = 16896;
        data[340] = 23552;
        data[341] = 0;
        data[342] = 16897;
        data[343] = 23552;
        data[344] = 514;
        data[345] = 17408;
        data[346] = 22019;
        data[347] = 18947;
        data[348] = 17920;
        data[349] = 17921;
        data[350] = 23040;
        data[351] = 17922;
        data[352] = 16898;
        data[353] = 23552;
        data[354] = 11780;
        data[355] = 41331;
        data[356] = 16897;
        data[357] = 23552;
        data[358] = 16896;
        data[359] = 23552;
        data[360] = 516;
        data[361] = 17408;
        data[362] = 16896;
        data[363] = 23552;
        data[364] = 518;
        data[365] = 17920;
        data[366] = 16898;
        data[367] = 23552;
        data[368] = 513;
        data[369] = 17922;
        data[370] = 33120;
        data[371] = 22019;
        data[372] = 18946;
        data[373] = 17920;
        data[374] = 17921;
        data[375] = 16896;
        data[376] = 23552;
        data[377] = 514;
        data[378] = 16384;
        data[379] = 23552;
        data[380] = 57824;
        data[381] = 14336;
        data[382] = 41369;
        data[383] = 49695;
        data[384] = 58344;
        data[385] = 15360;
        data[386] = 41368;
        data[387] = 57590;
        data[388] = 49695;
        data[389] = 3587;
        data[390] = 0;
        data[391] = 16384;
        data[392] = 23552;
        data[393] = 16896;
        data[394] = 23552;
        data[395] = 49499;
        data[396] = 16896;
        data[397] = 23552;
        data[398] = 516;
        data[399] = 16384;
        data[400] = 23552;
        data[401] = 3071;
        data[402] = 1546;
        data[403] = 16896;
        data[404] = 23552;
        data[405] = 514;
        data[406] = 17408;
        data[407] = 33176;
        data[408] = 33189;
        data[409] = 16896;
        data[410] = 23552;
        data[411] = 514;
        data[412] = 16384;
        data[413] = 23552;
        data[414] = 16897;
        data[415] = 23552;
        data[416] = 0;
        data[417] = 16896;
        data[418] = 23552;
        data[419] = 514;
        data[420] = 17408;
        data[421] = 22018;
        data[422] = 18946;
        data[423] = 17920;
        data[424] = 23040;
        data[425] = 17921;
        data[426] = 16897;
        data[427] = 23552;
        data[428] = 11780;
        data[429] = 41400;
        data[430] = 16897;
        data[431] = 23552;
        data[432] = 2566;
        data[433] = 514;
        data[434] = 49601;
        data[435] = 16897;
        data[436] = 23552;
        data[437] = 513;
        data[438] = 17921;
        data[439] = 33194;
        data[440] = 57611;
        data[441] = 16384;
        data[442] = 23552;
        data[443] = 16896;
        data[444] = 23552;
        data[445] = 0;
        data[446] = 57611;
        data[447] = 17408;
        data[448] = 22018;
        data[449] = 18945;
        data[450] = 17920;
        data[451] = 57611;
        data[452] = 16384;
        data[453] = 23552;
        data[454] = 57824;
        data[455] = 14336;
        data[456] = 41425;
        data[457] = 57611;
        data[458] = 16384;
        data[459] = 23552;
        data[460] = 57928;
        data[461] = 1024;
        data[462] = 57611;
        data[463] = 17408;
        data[464] = 33233;
        data[465] = 57611;
        data[466] = 16384;
        data[467] = 23552;
        data[468] = 65176;
        data[469] = 16896;
        data[470] = 23552;
        data[471] = 0;
        data[472] = 17408;
        data[473] = 57611;
        data[474] = 16384;
        data[475] = 23552;
        data[476] = 658;
        data[477] = 57611;
        data[478] = 17408;
        data[479] = 22017;
        data[480] = 18946;
        data[481] = 17920;
        data[482] = 17921;
        data[483] = 16896;
        data[484] = 23552;
        data[485] = 16897;
        data[486] = 23552;
        data[487] = 13312;
        data[488] = 41452;
        data[489] = 16896;
        data[490] = 23552;
        data[491] = 22018;
        data[492] = 16897;
        data[493] = 23552;
        data[494] = 22018;
        data[495] = 18946;
        data[496] = 17920;
        data[497] = 17921;
        data[498] = 16896;
        data[499] = 23552;
        data[500] = 16897;
        data[501] = 23552;
        data[502] = 11264;
        data[503] = 41467;
        data[504] = 16896;
        data[505] = 23552;
        data[506] = 22018;
        data[507] = 16897;
        data[508] = 23552;
        data[509] = 22018;
        data[510] = 18948;
        data[511] = 17920;
        data[512] = 17921;
        data[513] = 17922;
        data[514] = 16896;
        data[515] = 23552;
        data[516] = 16898;
        data[517] = 23552;
        data[518] = 0;
        data[519] = 17923;
        data[520] = 16896;
        data[521] = 23552;
        data[522] = 16899;
        data[523] = 23552;
        data[524] = 10240;
        data[525] = 41502;
        data[526] = 16896;
        data[527] = 23552;
        data[528] = 16384;
        data[529] = 23552;
        data[530] = 16897;
        data[531] = 23552;
        data[532] = 17408;
        data[533] = 16896;
        data[534] = 23552;
        data[535] = 513;
        data[536] = 17920;
        data[537] = 16897;
        data[538] = 23552;
        data[539] = 513;
        data[540] = 17921;
        data[541] = 33288;
        data[542] = 22020;
        data[543] = 57610;
        data[544] = 16384;
        data[545] = 23552;
        data[546] = 57610;
        data[547] = 16384;
        data[548] = 23552;
        data[549] = 6663;
        data[550] = 5120;
        data[551] = 57610;
        data[552] = 17408;
        data[553] = 57610;
        data[554] = 16384;
        data[555] = 23552;
        data[556] = 57610;
        data[557] = 16384;
        data[558] = 23552;
        data[559] = 7689;
        data[560] = 5120;
        data[561] = 57610;
        data[562] = 17408;
        data[563] = 57610;
        data[564] = 16384;
        data[565] = 23552;
        data[566] = 57610;
        data[567] = 16384;
        data[568] = 23552;
        data[569] = 6664;
        data[570] = 5120;
        data[571] = 57610;
        data[572] = 17408;
        data[573] = 57610;
        data[574] = 16384;
        data[575] = 23552;
        data[576] = 22016;

    end else begin
        // game data
        data[0] = 1;
        data[1] = 0;
        data[2] = 0;
        data[3] = 640;
        data[4] = 480;
        data[5] = 15139;
        data[6] = 1;
        data[7] = 207;
        data[8] = 0;
        data[9] = 225;
        data[10] = 480;
        data[11] = 13312;
        data[12] = 1;
        data[13] = 230;
        data[14] = 0;
        data[15] = 180;
        data[16] = 480;
        data[17] = 33808;
        data[18] = 1;
        data[19] = 245;
        data[20] = 0;
        data[21] = 150;
        data[22] = 480;
        data[23] = 40147;
        data[24] = 1;
        data[25] = 318;
        data[26] = 0;
        data[27] = 4;
        data[28] = 42;
        data[29] = 59196;
        data[30] = 1;
        data[31] = 318;
        data[32] = 146;
        data[33] = 4;
        data[34] = 42;
        data[35] = 59196;
        data[36] = 1;
        data[37] = 318;
        data[38] = 292;
        data[39] = 4;
        data[40] = 42;
        data[41] = 59196;
        data[42] = 1;
        data[43] = 318;
        data[44] = 438;
        data[45] = 4;
        data[46] = 42;
        data[47] = 59196;
        data[48] = 1;
        data[49] = 252;
        data[50] = 218;
        data[51] = 8;
        data[52] = 42;
        data[53] = 65120;
        data[54] = 0;
        data[55] = 32;
        data[56] = 0;
        data[57] = 8;
        data[58] = 42;
        data[59] = 59196;
        data[60] = 0;
        data[61] = 64;
        data[62] = 0;
        data[63] = 8;
        data[64] = 42;
        data[65] = 65120;
        data[66] = 0;
        data[67] = 96;
        data[68] = 0;
        data[69] = 8;
        data[70] = 42;
        data[71] = 59196;
        data[72] = 0;
        data[73] = 128;
        data[74] = 0;
        data[75] = 8;
        data[76] = 42;
        data[77] = 65120;
        data[78] = 1;
        data[79] = 60;
        data[80] = 140;
        data[81] = 80;
        data[82] = 200;
        data[83] = 20736;
        data[84] = 0;
        data[85] = -3;
        data[86] = -3;
        data[87] = 80;
        data[88] = 200;
        data[89] = 43552;
        data[90] = 0;
        data[91] = 35;
        data[92] = -3;
        data[93] = 4;
        data[94] = 200;
        data[95] = 53920;
        data[96] = 0;
        data[97] = 39;
        data[98] = -3;
        data[99] = 38;
        data[100] = 200;
        data[101] = 33152;
        data[102] = 1;
        data[103] = 500;
        data[104] = 140;
        data[105] = 80;
        data[106] = 200;
        data[107] = 20736;
        data[108] = 0;
        data[109] = -3;
        data[110] = -3;
        data[111] = 80;
        data[112] = 200;
        data[113] = 43552;
        data[114] = 0;
        data[115] = 35;
        data[116] = -3;
        data[117] = 4;
        data[118] = 200;
        data[119] = 53920;
        data[120] = 0;
        data[121] = 39;
        data[122] = -3;
        data[123] = 38;
        data[124] = 200;
        data[125] = 33152;
        data[126] = 1;
        data[127] = 348;
        data[128] = 350;
        data[129] = 24;
        data[130] = 9;
        data[131] = 0;
        data[132] = 0;
        data[133] = 0;
        data[134] = 32;
        data[135] = 24;
        data[136] = 9;
        data[137] = 0;
        data[138] = 0;
        data[139] = 2;
        data[140] = -8;
        data[141] = 20;
        data[142] = 56;
        data[143] = 63813;
        data[144] = 0;
        data[145] = 2;
        data[146] = -8;
        data[147] = 20;
        data[148] = 20;
        data[149] = 64170;
        data[150] = 0;
        data[151] = 2;
        data[152] = 7;
        data[153] = 20;
        data[154] = 6;
        data[155] = 64853;
        data[156] = 0;
        data[157] = 2;
        data[158] = 32;
        data[159] = 20;
        data[160] = 6;
        data[161] = 64853;
        data[162] = 1;
        data[163] = 348;
        data[164] = 100;
        data[165] = 24;
        data[166] = 9;
        data[167] = 0;
        data[168] = 0;
        data[169] = 0;
        data[170] = 32;
        data[171] = 24;
        data[172] = 9;
        data[173] = 0;
        data[174] = 0;
        data[175] = 2;
        data[176] = -8;
        data[177] = 20;
        data[178] = 54;
        data[179] = 1109;
        data[180] = 0;
        data[181] = 2;
        data[182] = 32;
        data[183] = 20;
        data[184] = 14;
        data[185] = 816;
        data[186] = 0;
        data[187] = 2;
        data[188] = 7;
        data[189] = 20;
        data[190] = 30;
        data[191] = 1370;
        data[192] = 0;
        data[193] = 4;
        data[194] = 14;
        data[195] = 16;
        data[196] = 18;
        data[197] = 816;
        data[198] = 1;
        data[199] = 260;
        data[200] = 0;
        data[201] = 40;
        data[202] = 128;
        data[203] = 816;
        data[204] = 0;
        data[205] = 10;
        data[206] = 128;
        data[207] = 20;
        data[208] = 4;
        data[209] = 0;
        data[210] = 0;
        data[211] = 0;
        data[212] = 155;
        data[213] = 40;
        data[214] = 9;
        data[215] = 0;
        data[216] = 0;
        data[217] = 2;
        data[218] = 132;
        data[219] = 36;
        data[220] = 40;
        data[221] = 1109;
        data[222] = 0;
        data[223] = 2;
        data[224] = 144;
        data[225] = 36;
        data[226] = 20;
        data[227] = 816;
        data[228] = 0;
        data[229] = 2;
        data[230] = 157;
        data[231] = 36;
        data[232] = 10;
        data[233] = 1370;
        data[234] = 0;
        data[235] = 5;
        data[236] = 157;
        data[237] = 30;
        data[238] = 4;
        data[239] = 816;
        data[240] = 0;
        data[241] = 2;
        data[242] = 166;
        data[243] = 36;
        data[244] = 6;
        data[245] = 1109;
        data[246] = 100;
        data[247] = 200;
        data[248] = 300;
        data[249] = 400;
        data[250] = 348;
        data[251] = 343;
        data[252] = 338;
        data[253] = 333;
        data[254] = 5;
        data[255] = 7;
        data[256] = 10;
        data[257] = 12;
        data[258] = 260;
        data[259] = 265;
        data[260] = 270;
        data[261] = 275;
        data[262] = 2;
        data[263] = 2;
        data[264] = 3;
        data[265] = 4;
        data[266] = 1;
        data[267] = 0;
        data[268] = 0;
        data[269] = 0;
        data[270] = 5;
        data[271] = 2;

    end
end


endmodule
