module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire [29:0] prom_inst_0_dout_w;
wire [29:0] prom_inst_1_dout_w;
wire [29:0] prom_inst_2_dout_w;
wire [29:0] prom_inst_3_dout_w;
wire [29:0] prom_inst_4_dout_w;
wire [29:0] prom_inst_5_dout_w;
wire [29:0] prom_inst_6_dout_w;
wire [29:0] prom_inst_7_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[29:0],dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 2;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hC2090CC824014F04B8C004A180D0000000008001001011004111041130411075;
defparam prom_inst_0.INIT_RAM_01 = 256'hD2A1092D02C0902C0901C0501939007C01F01407014052704000414440100830;
defparam prom_inst_0.INIT_RAM_02 = 256'h3C07C850180A0A468041A08C680E18082915122023C017F072005BC1C5108015;
defparam prom_inst_0.INIT_RAM_03 = 256'h04400704C03000C004080000000803C013C0130D1ECC072301C400557E0B01B1;
defparam prom_inst_0.INIT_RAM_04 = 256'h0300100C0B804038238910120C0000C00200003C02A20020090C040D0C040307;
defparam prom_inst_0.INIT_RAM_05 = 256'h030832001C020308908000098080304008228404C1200A30800C033030C40C10;
defparam prom_inst_0.INIT_RAM_06 = 256'h0043823CA16212A200A1061E1400842CD4280040CA000608001C108000100100;
defparam prom_inst_0.INIT_RAM_07 = 256'hC30810410010C109004AAA22F01305205019C1010401104800CC220440000340;
defparam prom_inst_0.INIT_RAM_08 = 256'h2C8232E8A12C8032E881AC8232E8812C823AE881ACAA6AAA48CCC40430420410;
defparam prom_inst_0.INIT_RAM_09 = 256'h00000000000000000000000000000000000000000000000000000000023AE8A1;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[29:0],dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 2;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h000010800000000002C000088000080010000000000011204112041110410313;
defparam prom_inst_1.INIT_RAM_01 = 256'h2010040100C02000030040000000003800C00C01000000300000100000000400;
defparam prom_inst_1.INIT_RAM_02 = 256'h1001083002080682002080A4201D0B0035012060000000100400044001011001;
defparam prom_inst_1.INIT_RAM_03 = 256'h0D014F0E812030840C1C0010010C1040C140C00841C10050401C400310040041;
defparam prom_inst_1.INIT_RAM_04 = 256'h0304A8001FC00100538F34F00010403103048404401910304F3C3C0B3C30024F;
defparam prom_inst_1.INIT_RAM_05 = 256'h0000910404120104406000420001110115564D30C330C3000404033030CC0C31;
defparam prom_inst_1.INIT_RAM_06 = 256'h04020F24B21002100230020A00100E40C8E800300E400300040000C000104404;
defparam prom_inst_1.INIT_RAM_07 = 256'hD0081681081D41D40C0797524B040C80CC3282000000000030C8310C43081101;
defparam prom_inst_1.INIT_RAM_08 = 256'h5B4B119430584F21A461594239B4B21A440984D31B51555D449AB10580400400;
defparam prom_inst_1.INIT_RAM_09 = 256'h00000000000000000000000000000000000000000000000000000000040584F3;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[29:0],dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 2;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h0000000000000000104000008000000000000000000011004110041100410001;
defparam prom_inst_2.INIT_RAM_01 = 256'h10300C0300802008010040100003003800F00802008000300200000000000400;
defparam prom_inst_2.INIT_RAM_02 = 256'h03003C30000B0E02C080B0102C100B0C10020000000000300000008002002002;
defparam prom_inst_2.INIT_RAM_03 = 256'h04C10707C11010440414000081001040B140B204408200A00004400303404004;
defparam prom_inst_2.INIT_RAM_04 = 256'h0104FC0009800024524924930C1000810104C00C00FC1010451C14051C140107;
defparam prom_inst_2.INIT_RAM_05 = 256'h030CF1000C320104407000074000010117FEC92C82208F30C000822010880421;
defparam prom_inst_2.INIT_RAM_06 = 256'h0441051010F109710840000400100C94ACC830F0C8C30E0C8C3433831030CC0E;
defparam prom_inst_2.INIT_RAM_07 = 256'hD00026026029029D000DBDF30C2006C0681343000000000020882308C20411C1;
defparam prom_inst_2.INIT_RAM_08 = 256'hB30C3F30D3F3092720B2F20913107171071F1020F01703D75047600980980940;
defparam prom_inst_2.INIT_RAM_09 = 256'h00000000000000000000000000000000000000000000000000000000030B00E3;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h0000004000000000104000000000000000000000000000000000000000000340;
defparam prom_inst_3.INIT_RAM_01 = 256'h0010000000000000000000000000000000000000000000300200080000000800;
defparam prom_inst_3.INIT_RAM_02 = 256'h0000043000070D01C34070901C14070C0401003000000020080000C031002001;
defparam prom_inst_3.INIT_RAM_03 = 256'h044107078110104404100000C100108020802004008200A0000800030080C00E;
defparam prom_inst_3.INIT_RAM_04 = 256'h010444000440001C60800400000000710104000000231010401C13041C10C107;
defparam prom_inst_3.INIT_RAM_05 = 256'h0000F0000C1300000030000DC00030001811010800000200000CC00010000401;
defparam prom_inst_3.INIT_RAM_06 = 256'h04010C34C3100710071000040000037C0C340000030000000008004000000000;
defparam prom_inst_3.INIT_RAM_07 = 256'hC0001001601C01C400044402662002C02C02C220000000001004000000001080;
defparam prom_inst_3.INIT_RAM_08 = 256'h92082D2092920B252092120921208292082D2092120D210140CFF00400580580;
defparam prom_inst_3.INIT_RAM_09 = 256'h000000000000000000000000000000000000000000000000000000000D3130A2;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[29:0],dout[9:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 2;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'h822AA808A822AA08880208A20AA2888A222888A222A8222082220822208283C8;
defparam prom_inst_4.INIT_RAM_01 = 256'hAA822AA822088220882208822AA820A0828220882208AAB2888AA28A88202022;
defparam prom_inst_4.INIT_RAM_02 = 256'h2A2AA4A2A924218908624218908624208628AA8222802A90AA00AA02B8AA8228;
defparam prom_inst_4.INIT_RAM_03 = 256'h06818705811010440418000841841A005A005A0628482A120A840AAAAA4ACAAD;
defparam prom_inst_4.INIT_RAM_04 = 256'h0106A8000A8000AC614514518628009101068008009910106A1C1A061C184187;
defparam prom_inst_4.INIT_RAM_05 = 256'h0106A280082A0208A0A0002A8000A28219CF8514411045104008411010440411;
defparam prom_inst_4.INIT_RAM_06 = 256'h04C18A24A242268226BA2A2E282AAE9AFACC10706CC10706C6141141B0104607;
defparam prom_inst_4.INIT_RAM_07 = 256'hE0208A08A08E08E02AA0E0EBFFBE03A0380BCB20208202AA304C1304C18C1363;
defparam prom_inst_4.INIT_RAM_08 = 256'h4289282892828A2828A2428A2828A2428A2828A2828C28787AFEE82282282242;
defparam prom_inst_4.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000089282892;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[29:0],dout[11:10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 2;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h48856022118858E20428E21121884E213884E213886204682047820468200C05;
defparam prom_inst_5.INIT_RAM_01 = 256'h5608856188621886218862188561861618588621886216282061812121888388;
defparam prom_inst_5.INIT_RAM_02 = 256'h4A80A1A8608080602018080602018082008456088849849A252612E8B4560884;
defparam prom_inst_5.INIT_RAM_03 = 256'h80201280A0420810820182022022031803180180491882066091618A0A126024;
defparam prom_inst_5.INIT_RAM_04 = 256'h208001820018200114104104514520042080120120004208004A00804A022012;
defparam prom_inst_5.INIT_RAM_05 = 256'h2080045202302081080608001820042044CF5041204810481202204208108204;
defparam prom_inst_5.INIT_RAM_06 = 256'h81E01D71D70283428344858286058000000E080800E080801142042002081080;
defparam prom_inst_5.INIT_RAM_07 = 256'h88860560560560508580D0D0000E80E80E00208886088858781E0781E01E0707;
defparam prom_inst_5.INIT_RAM_08 = 256'h035C7435C7435D7435D7035D7035D7035D7435D7435034343433318158158118;
defparam prom_inst_5.INIT_RAM_09 = 256'h000000000000000000000000000000000000000000000000000000001C7035C7;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[29:0],dout[13:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 2;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'h044004110044011100B411001014151054415105440522549225492254924424;
defparam prom_inst_6.INIT_RAM_01 = 256'h50444404441104411044110440044111044441104411004452D0101010444A44;
defparam prom_inst_6.INIT_RAM_02 = 256'h97457A7404404A9012A404A9012A40412B405044440045711C0115C470504440;
defparam prom_inst_6.INIT_RAM_03 = 256'h4AD2084AD2212488492A4927927926048604844997A745E9D17A901757A5D15E;
defparam prom_inst_6.INIT_RAM_04 = 256'h12490A4920A49240928A28A249249282124909209288212490212B48212B9208;
defparam prom_inst_6.INIT_RAM_05 = 256'h524902492936D24884A92490A492421224CF4A2092248824892B922124884922;
defparam prom_inst_6.INIT_RAM_06 = 256'h48D24D38D3804B404B40404B41211001010D24A490D24A49092122126D24884A;
defparam prom_inst_6.INIT_RAM_07 = 256'h04410510510510524412D2D4004C48C48D2412E441044401348D2348D24D2313;
defparam prom_inst_6.INIT_RAM_08 = 256'h8B4E34B4E34B4D34B4D38B4D38B4D38B4D34B4D34B40B4B4B533344144144184;
defparam prom_inst_6.INIT_RAM_09 = 256'h000000000000000000000000000000000000000000000000000000004E38B4E3;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[29:0],dout[15:14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 2;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'h455554D5505555156785155DD55541550554155055557705D7705D7705D767E7;
defparam prom_inst_7.INIT_RAM_01 = 256'h5575555555555555555555555555515545555555555555455615591515555855;
defparam prom_inst_7.INIT_RAM_02 = 256'h03543835575B5E16D785B5E16D785B5D78575575554054314D0150C537557557;
defparam prom_inst_7.INIT_RAM_03 = 256'h5E179C5E177175DC5D785D74D74D74C5F4C5F45DD38354E0D538D5534380D50E;
defparam prom_inst_7.INIT_RAM_04 = 256'h175DB85D7B85D76DD7DF7DF75D75D7B7175D9D79D7BB7175DA71785E7178D79C;
defparam prom_inst_7.INIT_RAM_05 = 256'h175DA75D7976175DC5E175DB85D7671777FF5F7DD775DF75DD78D77175DC5D77;
defparam prom_inst_7.INIT_RAM_06 = 256'h5DD75D7DD7F05F705F64545855755FFDFDBD75E5DBD75E5D9D7D77D76175DC5E;
defparam prom_inst_7.INIT_RAM_07 = 256'h055575575575575F555FDFD7FF7C5FC5FD76D6355545555575DD775DD75D77D7;
defparam prom_inst_7.INIT_RAM_08 = 256'hFF5F77F5F77F5D77F5D7FF5D7FF5D7FF5D77F5D77F7FF7F7F5FFF55D55D55DD5;
defparam prom_inst_7.INIT_RAM_09 = 256'h000000000000000000000000000000000000000000000000000000005F7FF5F7;

endmodule //Gowin_pROM
