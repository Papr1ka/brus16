/*
    1*READ 1*WRITE sync memory
    intended to be implemented as block ram
    sync read, sync write
*/

module bsram
#(
    parameter WIDTH = 13,
    parameter SIZE = 8192,
    parameter LOAD_PROGRAM = 1
)
(
    input wire clk,

    // read
    input wire [WIDTH-1:0] mem_dout_addr,
    output reg [15:0] mem_dout,
    
    // write
    input wire we,
    input wire [WIDTH-1:0] mem_din_addr,
    input wire [15:0] mem_din
);

reg [15:0] data [SIZE-1:0];

always_ff @(posedge clk) begin
    if (we) begin
        data[mem_din_addr] <= mem_din;
    end
    mem_dout <= data[mem_dout_addr];
end

initial begin
    for (integer i = 0; i < SIZE; i = i + 1) begin
        data[i] = 16'b0;
    end
    if (LOAD_PROGRAM) begin
        // game program
        data[0] = 65136;
        data[1] = 19456;
        data[2] = 49161;
        data[3] = 23041;
        data[4] = 40968;
        data[5] = 49166;
        data[6] = 25600;
        data[7] = 32771;
        data[8] = 22016;
        data[9] = 23286;
        data[10] = 65152;
        data[11] = 57344;
        data[12] = 49858;
        data[13] = 22016;
        data[14] = 49397;
        data[15] = 49172;
        data[16] = 49236;
        data[17] = 49581;
        data[18] = 49294;
        data[19] = 22016;
        data[20] = 65136;
        data[21] = 16384;
        data[22] = 23552;
        data[23] = 40991;
        data[24] = 57597;
        data[25] = 16384;
        data[26] = 23552;
        data[27] = 522;
        data[28] = 57597;
        data[29] = 17408;
        data[30] = 32799;
        data[31] = 65137;
        data[32] = 16384;
        data[33] = 23552;
        data[34] = 41005;
        data[35] = 57597;
        data[36] = 16384;
        data[37] = 23552;
        data[38] = 1556;
        data[39] = 57597;
        data[40] = 17408;
        data[41] = 23040;
        data[42] = 57596;
        data[43] = 17408;
        data[44] = 32813;
        data[45] = 65138;
        data[46] = 16384;
        data[47] = 23552;
        data[48] = 41019;
        data[49] = 57597;
        data[50] = 16384;
        data[51] = 23552;
        data[52] = 14948;
        data[53] = 41018;
        data[54] = 23522;
        data[55] = 57596;
        data[56] = 17408;
        data[57] = 32826;
        data[58] = 32827;
        data[59] = 65139;
        data[60] = 16384;
        data[61] = 23552;
        data[62] = 41033;
        data[63] = 57597;
        data[64] = 16384;
        data[65] = 23552;
        data[66] = 14948;
        data[67] = 41032;
        data[68] = 23070;
        data[69] = 57596;
        data[70] = 17408;
        data[71] = 32840;
        data[72] = 32841;
        data[73] = 57597;
        data[74] = 16384;
        data[75] = 23552;
        data[76] = 1539;
        data[77] = 23040;
        data[78] = 49828;
        data[79] = 59344;
        data[80] = 49843;
        data[81] = 57597;
        data[82] = 17408;
        data[83] = 22016;
        data[84] = 18946;
        data[85] = 23041;
        data[86] = 59344;
        data[87] = 57597;
        data[88] = 16384;
        data[89] = 23552;
        data[90] = 1024;
        data[91] = 7689;
        data[92] = 0;
        data[93] = 17920;
        data[94] = 57596;
        data[95] = 16384;
        data[96] = 23552;
        data[97] = 13824;
        data[98] = 41070;
        data[99] = 57596;
        data[100] = 16384;
        data[101] = 23552;
        data[102] = 16896;
        data[103] = 23552;
        data[104] = 1024;
        data[105] = 23040;
        data[106] = 49828;
        data[107] = 57596;
        data[108] = 17408;
        data[109] = 32894;
        data[110] = 57596;
        data[111] = 16384;
        data[112] = 23552;
        data[113] = 11776;
        data[114] = 41086;
        data[115] = 57596;
        data[116] = 16384;
        data[117] = 23552;
        data[118] = 16896;
        data[119] = 23552;
        data[120] = 0;
        data[121] = 23040;
        data[122] = 49843;
        data[123] = 57596;
        data[124] = 17408;
        data[125] = 32894;
        data[126] = 65279;
        data[127] = 16384;
        data[128] = 23552;
        data[129] = 17921;
        data[130] = 16897;
        data[131] = 23552;
        data[132] = 57596;
        data[133] = 16384;
        data[134] = 23552;
        data[135] = 516;
        data[136] = 23043;
        data[137] = 8192;
        data[138] = 0;
        data[139] = 65279;
        data[140] = 17408;
        data[141] = 22018;
        data[142] = 58344;
        data[143] = 57602;
        data[144] = 57598;
        data[145] = 23472;
        data[146] = 58324;
        data[147] = 23294;
        data[148] = 6664;
        data[149] = 4620;
        data[150] = 65314;
        data[151] = 49315;
        data[152] = 57844;
        data[153] = 57611;
        data[154] = 57607;
        data[155] = 23352;
        data[156] = 57824;
        data[157] = 23294;
        data[158] = 6664;
        data[159] = 4620;
        data[160] = 65350;
        data[161] = 49315;
        data[162] = 22016;
        data[163] = 18951;
        data[164] = 17920;
        data[165] = 17921;
        data[166] = 17922;
        data[167] = 17923;
        data[168] = 17924;
        data[169] = 17925;
        data[170] = 17926;
        data[171] = 16896;
        data[172] = 23552;
        data[173] = 514;
        data[174] = 16384;
        data[175] = 23552;
        data[176] = 16898;
        data[177] = 23552;
        data[178] = 14336;
        data[179] = 16896;
        data[180] = 23552;
        data[181] = 514;
        data[182] = 16384;
        data[183] = 23552;
        data[184] = 16897;
        data[185] = 23552;
        data[186] = 12288;
        data[187] = 4096;
        data[188] = 41185;
        data[189] = 49891;
        data[190] = 16902;
        data[191] = 23552;
        data[192] = 15360;
        data[193] = 41184;
        data[194] = 16900;
        data[195] = 23552;
        data[196] = 49891;
        data[197] = 3587;
        data[198] = 0;
        data[199] = 16384;
        data[200] = 23552;
        data[201] = 16896;
        data[202] = 23552;
        data[203] = 513;
        data[204] = 17408;
        data[205] = 16899;
        data[206] = 23552;
        data[207] = 16896;
        data[208] = 23552;
        data[209] = 514;
        data[210] = 17408;
        data[211] = 16901;
        data[212] = 23552;
        data[213] = 23041;
        data[214] = 49891;
        data[215] = 3587;
        data[216] = 0;
        data[217] = 0;
        data[218] = 16384;
        data[219] = 23552;
        data[220] = 16901;
        data[221] = 23552;
        data[222] = 17408;
        data[223] = 32992;
        data[224] = 33012;
        data[225] = 16896;
        data[226] = 23552;
        data[227] = 514;
        data[228] = 16384;
        data[229] = 23552;
        data[230] = 16901;
        data[231] = 23552;
        data[232] = 16384;
        data[233] = 23552;
        data[234] = 57597;
        data[235] = 16384;
        data[236] = 23552;
        data[237] = 7687;
        data[238] = 0;
        data[239] = 0;
        data[240] = 16896;
        data[241] = 23552;
        data[242] = 514;
        data[243] = 17408;
        data[244] = 22023;
        data[245] = 18959;
        data[246] = 65278;
        data[247] = 17920;
        data[248] = 16896;
        data[249] = 23552;
        data[250] = 513;
        data[251] = 16384;
        data[252] = 23552;
        data[253] = 514;
        data[254] = 17921;
        data[255] = 16896;
        data[256] = 23552;
        data[257] = 514;
        data[258] = 16384;
        data[259] = 23552;
        data[260] = 1016;
        data[261] = 17922;
        data[262] = 16897;
        data[263] = 23552;
        data[264] = 532;
        data[265] = 17923;
        data[266] = 16898;
        data[267] = 23552;
        data[268] = 568;
        data[269] = 17924;
        data[270] = 16897;
        data[271] = 23552;
        data[272] = 12006;
        data[273] = 16899;
        data[274] = 23552;
        data[275] = 57754;
        data[276] = 13312;
        data[277] = 4096;
        data[278] = 41241;
        data[279] = 49519;
        data[280] = 33049;
        data[281] = 65314;
        data[282] = 17925;
        data[283] = 16901;
        data[284] = 23552;
        data[285] = 513;
        data[286] = 16384;
        data[287] = 23552;
        data[288] = 17926;
        data[289] = 16901;
        data[290] = 23552;
        data[291] = 514;
        data[292] = 16384;
        data[293] = 23552;
        data[294] = 1016;
        data[295] = 17927;
        data[296] = 16902;
        data[297] = 23552;
        data[298] = 536;
        data[299] = 17928;
        data[300] = 16903;
        data[301] = 23552;
        data[302] = 566;
        data[303] = 17929;
        data[304] = 16905;
        data[305] = 23552;
        data[306] = 16904;
        data[307] = 23552;
        data[308] = 16903;
        data[309] = 23552;
        data[310] = 16902;
        data[311] = 23552;
        data[312] = 16900;
        data[313] = 23552;
        data[314] = 16899;
        data[315] = 23552;
        data[316] = 16898;
        data[317] = 23552;
        data[318] = 16897;
        data[319] = 23552;
        data[320] = 49785;
        data[321] = 41284;
        data[322] = 49519;
        data[323] = 33092;
        data[324] = 65350;
        data[325] = 17930;
        data[326] = 16906;
        data[327] = 23552;
        data[328] = 513;
        data[329] = 16384;
        data[330] = 23552;
        data[331] = 17931;
        data[332] = 16906;
        data[333] = 23552;
        data[334] = 514;
        data[335] = 16384;
        data[336] = 23552;
        data[337] = 17932;
        data[338] = 16907;
        data[339] = 23552;
        data[340] = 552;
        data[341] = 17933;
        data[342] = 16908;
        data[343] = 23552;
        data[344] = 684;
        data[345] = 17934;
        data[346] = 16910;
        data[347] = 23552;
        data[348] = 16909;
        data[349] = 23552;
        data[350] = 16908;
        data[351] = 23552;
        data[352] = 16907;
        data[353] = 23552;
        data[354] = 16900;
        data[355] = 23552;
        data[356] = 16899;
        data[357] = 23552;
        data[358] = 16898;
        data[359] = 23552;
        data[360] = 16897;
        data[361] = 23552;
        data[362] = 49785;
        data[363] = 41326;
        data[364] = 49519;
        data[365] = 33134;
        data[366] = 22031;
        data[367] = 18948;
        data[368] = 65278;
        data[369] = 17920;
        data[370] = 16896;
        data[371] = 23552;
        data[372] = 514;
        data[373] = 16384;
        data[374] = 23552;
        data[375] = 17921;
        data[376] = 23040;
        data[377] = 17922;
        data[378] = 16898;
        data[379] = 23552;
        data[380] = 11781;
        data[381] = 41384;
        data[382] = 23040;
        data[383] = 17923;
        data[384] = 16897;
        data[385] = 23552;
        data[386] = 16896;
        data[387] = 23552;
        data[388] = 514;
        data[389] = 17408;
        data[390] = 16899;
        data[391] = 23552;
        data[392] = 11791;
        data[393] = 41360;
        data[394] = 25600;
        data[395] = 16899;
        data[396] = 23552;
        data[397] = 513;
        data[398] = 17923;
        data[399] = 33158;
        data[400] = 23040;
        data[401] = 17923;
        data[402] = 23292;
        data[403] = 6664;
        data[404] = 4632;
        data[405] = 16896;
        data[406] = 23552;
        data[407] = 514;
        data[408] = 17408;
        data[409] = 16899;
        data[410] = 23552;
        data[411] = 11806;
        data[412] = 41379;
        data[413] = 25600;
        data[414] = 16899;
        data[415] = 23552;
        data[416] = 513;
        data[417] = 17923;
        data[418] = 33177;
        data[419] = 16898;
        data[420] = 23552;
        data[421] = 513;
        data[422] = 17922;
        data[423] = 33146;
        data[424] = 23041;
        data[425] = 41388;
        data[426] = 25600;
        data[427] = 33192;
        data[428] = 22020;
        data[429] = 18945;
        data[430] = 57597;
        data[431] = 16384;
        data[432] = 23552;
        data[433] = 7687;
        data[434] = 17920;
        data[435] = 16896;
        data[436] = 23552;
        data[437] = 49727;
        data[438] = 16896;
        data[439] = 23552;
        data[440] = 49602;
        data[441] = 16896;
        data[442] = 23552;
        data[443] = 65230;
        data[444] = 49677;
        data[445] = 16896;
        data[446] = 23552;
        data[447] = 65254;
        data[448] = 49677;
        data[449] = 22017;
        data[450] = 18947;
        data[451] = 17920;
        data[452] = 65200;
        data[453] = 17921;
        data[454] = 65176;
        data[455] = 17922;
        data[456] = 16897;
        data[457] = 23552;
        data[458] = 514;
        data[459] = 16384;
        data[460] = 23552;
        data[461] = 57824;
        data[462] = 14336;
        data[463] = 49891;
        data[464] = 58344;
        data[465] = 15360;
        data[466] = 3072;
        data[467] = 41447;
        data[468] = 16898;
        data[469] = 23552;
        data[470] = 514;
        data[471] = 16384;
        data[472] = 23552;
        data[473] = 11776;
        data[474] = 41446;
        data[475] = 16898;
        data[476] = 23552;
        data[477] = 514;
        data[478] = 16384;
        data[479] = 23552;
        data[480] = 1609;
        data[481] = 16897;
        data[482] = 23552;
        data[483] = 514;
        data[484] = 17408;
        data[485] = 33254;
        data[486] = 33255;
        data[487] = 16897;
        data[488] = 23552;
        data[489] = 514;
        data[490] = 16384;
        data[491] = 23552;
        data[492] = 16896;
        data[493] = 23552;
        data[494] = 0;
        data[495] = 16897;
        data[496] = 23552;
        data[497] = 514;
        data[498] = 17408;
        data[499] = 22019;
        data[500] = 18947;
        data[501] = 17920;
        data[502] = 17921;
        data[503] = 23040;
        data[504] = 17922;
        data[505] = 16898;
        data[506] = 23552;
        data[507] = 11780;
        data[508] = 41484;
        data[509] = 16897;
        data[510] = 23552;
        data[511] = 16896;
        data[512] = 23552;
        data[513] = 516;
        data[514] = 17408;
        data[515] = 16896;
        data[516] = 23552;
        data[517] = 518;
        data[518] = 17920;
        data[519] = 16898;
        data[520] = 23552;
        data[521] = 513;
        data[522] = 17922;
        data[523] = 33273;
        data[524] = 22019;
        data[525] = 18946;
        data[526] = 17920;
        data[527] = 17921;
        data[528] = 16896;
        data[529] = 23552;
        data[530] = 514;
        data[531] = 16384;
        data[532] = 23552;
        data[533] = 57824;
        data[534] = 14336;
        data[535] = 41522;
        data[536] = 49891;
        data[537] = 58344;
        data[538] = 15360;
        data[539] = 41521;
        data[540] = 57590;
        data[541] = 49891;
        data[542] = 3587;
        data[543] = 0;
        data[544] = 16384;
        data[545] = 23552;
        data[546] = 16896;
        data[547] = 23552;
        data[548] = 49652;
        data[549] = 16896;
        data[550] = 23552;
        data[551] = 516;
        data[552] = 16384;
        data[553] = 23552;
        data[554] = 3071;
        data[555] = 1546;
        data[556] = 16896;
        data[557] = 23552;
        data[558] = 514;
        data[559] = 17408;
        data[560] = 33329;
        data[561] = 33342;
        data[562] = 16896;
        data[563] = 23552;
        data[564] = 514;
        data[565] = 16384;
        data[566] = 23552;
        data[567] = 16897;
        data[568] = 23552;
        data[569] = 0;
        data[570] = 16896;
        data[571] = 23552;
        data[572] = 514;
        data[573] = 17408;
        data[574] = 22018;
        data[575] = 18946;
        data[576] = 17920;
        data[577] = 23040;
        data[578] = 17921;
        data[579] = 16897;
        data[580] = 23552;
        data[581] = 11780;
        data[582] = 41553;
        data[583] = 16897;
        data[584] = 23552;
        data[585] = 2566;
        data[586] = 514;
        data[587] = 49754;
        data[588] = 16897;
        data[589] = 23552;
        data[590] = 513;
        data[591] = 17921;
        data[592] = 33347;
        data[593] = 57595;
        data[594] = 16384;
        data[595] = 23552;
        data[596] = 16896;
        data[597] = 23552;
        data[598] = 0;
        data[599] = 57595;
        data[600] = 17408;
        data[601] = 22018;
        data[602] = 18945;
        data[603] = 17920;
        data[604] = 57595;
        data[605] = 16384;
        data[606] = 23552;
        data[607] = 57824;
        data[608] = 14336;
        data[609] = 41578;
        data[610] = 57595;
        data[611] = 16384;
        data[612] = 23552;
        data[613] = 57928;
        data[614] = 1024;
        data[615] = 57595;
        data[616] = 17408;
        data[617] = 33386;
        data[618] = 57595;
        data[619] = 16384;
        data[620] = 23552;
        data[621] = 65176;
        data[622] = 16896;
        data[623] = 23552;
        data[624] = 0;
        data[625] = 17408;
        data[626] = 57595;
        data[627] = 16384;
        data[628] = 23552;
        data[629] = 658;
        data[630] = 57595;
        data[631] = 17408;
        data[632] = 22017;
        data[633] = 18952;
        data[634] = 17920;
        data[635] = 17921;
        data[636] = 17922;
        data[637] = 17923;
        data[638] = 17924;
        data[639] = 17925;
        data[640] = 17926;
        data[641] = 17927;
        data[642] = 16898;
        data[643] = 23552;
        data[644] = 16900;
        data[645] = 23552;
        data[646] = 11264;
        data[647] = 41610;
        data[648] = 23040;
        data[649] = 22024;
        data[650] = 16896;
        data[651] = 23552;
        data[652] = 16902;
        data[653] = 23552;
        data[654] = 13312;
        data[655] = 41618;
        data[656] = 23040;
        data[657] = 22024;
        data[658] = 16899;
        data[659] = 23552;
        data[660] = 16901;
        data[661] = 23552;
        data[662] = 11264;
        data[663] = 41626;
        data[664] = 23040;
        data[665] = 22024;
        data[666] = 16897;
        data[667] = 23552;
        data[668] = 16903;
        data[669] = 23552;
        data[670] = 13312;
        data[671] = 41634;
        data[672] = 23040;
        data[673] = 22024;
        data[674] = 23041;
        data[675] = 22024;
        data[676] = 18946;
        data[677] = 17920;
        data[678] = 17921;
        data[679] = 16896;
        data[680] = 23552;
        data[681] = 16897;
        data[682] = 23552;
        data[683] = 13312;
        data[684] = 41648;
        data[685] = 16896;
        data[686] = 23552;
        data[687] = 22018;
        data[688] = 16897;
        data[689] = 23552;
        data[690] = 22018;
        data[691] = 18946;
        data[692] = 17920;
        data[693] = 17921;
        data[694] = 16896;
        data[695] = 23552;
        data[696] = 16897;
        data[697] = 23552;
        data[698] = 11264;
        data[699] = 41663;
        data[700] = 16896;
        data[701] = 23552;
        data[702] = 22018;
        data[703] = 16897;
        data[704] = 23552;
        data[705] = 22018;
        data[706] = 18948;
        data[707] = 17920;
        data[708] = 17921;
        data[709] = 17922;
        data[710] = 16896;
        data[711] = 23552;
        data[712] = 16898;
        data[713] = 23552;
        data[714] = 0;
        data[715] = 17923;
        data[716] = 16896;
        data[717] = 23552;
        data[718] = 16899;
        data[719] = 23552;
        data[720] = 10240;
        data[721] = 41698;
        data[722] = 16896;
        data[723] = 23552;
        data[724] = 16384;
        data[725] = 23552;
        data[726] = 16897;
        data[727] = 23552;
        data[728] = 17408;
        data[729] = 16896;
        data[730] = 23552;
        data[731] = 513;
        data[732] = 17920;
        data[733] = 16897;
        data[734] = 23552;
        data[735] = 513;
        data[736] = 17921;
        data[737] = 33484;
        data[738] = 22020;
        data[739] = 57594;
        data[740] = 16384;
        data[741] = 23552;
        data[742] = 57594;
        data[743] = 16384;
        data[744] = 23552;
        data[745] = 6663;
        data[746] = 5120;
        data[747] = 57594;
        data[748] = 17408;
        data[749] = 57594;
        data[750] = 16384;
        data[751] = 23552;
        data[752] = 57594;
        data[753] = 16384;
        data[754] = 23552;
        data[755] = 7689;
        data[756] = 5120;
        data[757] = 57594;
        data[758] = 17408;
        data[759] = 57594;
        data[760] = 16384;
        data[761] = 23552;
        data[762] = 57594;
        data[763] = 16384;
        data[764] = 23552;
        data[765] = 6664;
        data[766] = 5120;
        data[767] = 57594;
        data[768] = 17408;
        data[769] = 57594;
        data[770] = 16384;
        data[771] = 23552;
        data[772] = 22016;

    end else begin
        // game data
		data[0] = 1;
        data[1] = 0;
        data[2] = 0;
        data[3] = 640;
        data[4] = 480;
        data[5] = 15139;
        data[6] = 1;
        data[7] = 207;
        data[8] = 0;
        data[9] = 225;
        data[10] = 480;
        data[11] = 13312;
        data[12] = 1;
        data[13] = 230;
        data[14] = 0;
        data[15] = 180;
        data[16] = 480;
        data[17] = 33808;
        data[18] = 1;
        data[19] = 245;
        data[20] = 0;
        data[21] = 150;
        data[22] = 480;
        data[23] = 40147;
        data[24] = 1;
        data[25] = 318;
        data[26] = 0;
        data[27] = 4;
        data[28] = 42;
        data[29] = 59196;
        data[30] = 1;
        data[31] = 318;
        data[32] = 146;
        data[33] = 4;
        data[34] = 42;
        data[35] = 59196;
        data[36] = 1;
        data[37] = 318;
        data[38] = 292;
        data[39] = 4;
        data[40] = 42;
        data[41] = 59196;
        data[42] = 1;
        data[43] = 318;
        data[44] = 438;
        data[45] = 4;
        data[46] = 42;
        data[47] = 59196;
        data[48] = 1;
        data[49] = 252;
        data[50] = 218;
        data[51] = 8;
        data[52] = 42;
        data[53] = 65120;
        data[54] = 0;
        data[55] = 32;
        data[56] = 0;
        data[57] = 8;
        data[58] = 42;
        data[59] = 59196;
        data[60] = 0;
        data[61] = 64;
        data[62] = 0;
        data[63] = 8;
        data[64] = 42;
        data[65] = 65120;
        data[66] = 0;
        data[67] = 96;
        data[68] = 0;
        data[69] = 8;
        data[70] = 42;
        data[71] = 59196;
        data[72] = 0;
        data[73] = 128;
        data[74] = 0;
        data[75] = 8;
        data[76] = 42;
        data[77] = 65120;
        data[78] = 1;
        data[79] = 60;
        data[80] = 140;
        data[81] = 80;
        data[82] = 200;
        data[83] = 20736;
        data[84] = 0;
        data[85] = 65533;
        data[86] = 65533;
        data[87] = 80;
        data[88] = 200;
        data[89] = 43552;
        data[90] = 0;
        data[91] = 35;
        data[92] = 65533;
        data[93] = 4;
        data[94] = 200;
        data[95] = 53920;
        data[96] = 0;
        data[97] = 39;
        data[98] = 65533;
        data[99] = 38;
        data[100] = 200;
        data[101] = 33152;
        data[102] = 1;
        data[103] = 500;
        data[104] = 140;
        data[105] = 80;
        data[106] = 200;
        data[107] = 20736;
        data[108] = 0;
        data[109] = 65533;
        data[110] = 65533;
        data[111] = 80;
        data[112] = 200;
        data[113] = 43552;
        data[114] = 0;
        data[115] = 35;
        data[116] = 65533;
        data[117] = 4;
        data[118] = 200;
        data[119] = 53920;
        data[120] = 0;
        data[121] = 39;
        data[122] = 65533;
        data[123] = 38;
        data[124] = 200;
        data[125] = 33152;
        data[126] = 1;
        data[127] = 348;
        data[128] = 350;
        data[129] = 24;
        data[130] = 9;
        data[131] = 0;
        data[132] = 0;
        data[133] = 0;
        data[134] = 32;
        data[135] = 24;
        data[136] = 9;
        data[137] = 0;
        data[138] = 0;
        data[139] = 2;
        data[140] = 65528;
        data[141] = 20;
        data[142] = 56;
        data[143] = 63813;
        data[144] = 0;
        data[145] = 2;
        data[146] = 65528;
        data[147] = 20;
        data[148] = 20;
        data[149] = 64170;
        data[150] = 0;
        data[151] = 2;
        data[152] = 7;
        data[153] = 20;
        data[154] = 6;
        data[155] = 64853;
        data[156] = 0;
        data[157] = 2;
        data[158] = 32;
        data[159] = 20;
        data[160] = 6;
        data[161] = 64853;
        data[162] = 1;
        data[163] = 348;
        data[164] = 100;
        data[165] = 24;
        data[166] = 9;
        data[167] = 0;
        data[168] = 0;
        data[169] = 0;
        data[170] = 32;
        data[171] = 24;
        data[172] = 9;
        data[173] = 0;
        data[174] = 0;
        data[175] = 2;
        data[176] = 65528;
        data[177] = 20;
        data[178] = 54;
        data[179] = 1109;
        data[180] = 0;
        data[181] = 2;
        data[182] = 32;
        data[183] = 20;
        data[184] = 14;
        data[185] = 816;
        data[186] = 0;
        data[187] = 2;
        data[188] = 7;
        data[189] = 20;
        data[190] = 30;
        data[191] = 1370;
        data[192] = 0;
        data[193] = 4;
        data[194] = 14;
        data[195] = 16;
        data[196] = 18;
        data[197] = 816;
        data[198] = 1;
        data[199] = 260;
        data[200] = 200;
        data[201] = 40;
        data[202] = 128;
        data[203] = 816;
        data[204] = 0;
        data[205] = 10;
        data[206] = 128;
        data[207] = 20;
        data[208] = 4;
        data[209] = 0;
        data[210] = 0;
        data[211] = 0;
        data[212] = 155;
        data[213] = 40;
        data[214] = 9;
        data[215] = 0;
        data[216] = 0;
        data[217] = 2;
        data[218] = 132;
        data[219] = 36;
        data[220] = 40;
        data[221] = 1109;
        data[222] = 0;
        data[223] = 2;
        data[224] = 144;
        data[225] = 36;
        data[226] = 20;
        data[227] = 816;
        data[228] = 0;
        data[229] = 2;
        data[230] = 157;
        data[231] = 36;
        data[232] = 10;
        data[233] = 1370;
        data[234] = 0;
        data[235] = 5;
        data[236] = 157;
        data[237] = 30;
        data[238] = 4;
        data[239] = 816;
        data[240] = 0;
        data[241] = 2;
        data[242] = 166;
        data[243] = 36;
        data[244] = 6;
        data[245] = 1109;
        data[246] = 100;
        data[247] = 200;
        data[248] = 300;
        data[249] = 400;
        data[250] = 1;
        data[251] = 0;
        data[252] = 0;
        data[253] = 0;
        data[254] = 348;
        data[255] = 368;
        data[256] = 338;
        data[257] = 328;
        data[258] = 65531;
        data[259] = 65531;
        data[260] = 65529;
        data[261] = 65526;
        data[262] = 65524;
        data[263] = 260;
        data[264] = 245;
        data[265] = 270;
        data[266] = 280;
        data[267] = 2;
        data[268] = 2;
        data[269] = 2;
        data[270] = 3;
        data[271] = 4;
    end
end


endmodule
