//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Sun Oct 26 14:24:20 2025

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire [29:0] prom_inst_0_dout_w;
wire [29:0] prom_inst_1_dout_w;
wire [29:0] prom_inst_2_dout_w;
wire [29:0] prom_inst_3_dout_w;
wire [29:0] prom_inst_4_dout_w;
wire [29:0] prom_inst_5_dout_w;
wire [29:0] prom_inst_6_dout_w;
wire [29:0] prom_inst_7_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[29:0],dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 2;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h3820002008300020004046063305020050F82807090040507181C0100108C850;
defparam prom_inst_0.INIT_RAM_01 = 256'h06040BC803040420F0403912031003830A00420082093932820F2820A2330014;
defparam prom_inst_0.INIT_RAM_02 = 256'h734A10808D9048C0C04A010C08B04ABB048C08C058C0B02181162023840B0602;
defparam prom_inst_0.INIT_RAM_03 = 256'h01C284F210021921422408A02008610D20204203053359234CA320031D33CC80;
defparam prom_inst_0.INIT_RAM_04 = 256'h93904E0C000D300D00C63003945A101429082C00C00E80900808010812C92200;
defparam prom_inst_0.INIT_RAM_05 = 256'h2008221082230823511004010C3082421820412860C1048410C4104C1080100B;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000002;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[29:0],dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 2;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h3CC000F03CC000F03080C00C000E8F90E028C90E0330D0F03383C03D50040E20;
defparam prom_inst_1.INIT_RAM_01 = 256'h00000F40010C0400304000100000000704000000000540107B2643B4C8304300;
defparam prom_inst_1.INIT_RAM_02 = 256'h01400000DFF800048CCFCF8B00A00A4C80004448A46858014014B82041804080;
defparam prom_inst_1.INIT_RAM_03 = 256'h00900000000005008004001080000800D0F003010C522008003000AC1003C000;
defparam prom_inst_1.INIT_RAM_04 = 256'h54020808020A220A008020020021010003C02C10000072300000000000200101;
defparam prom_inst_1.INIT_RAM_05 = 256'h220822208221082600000000000000040030000000C000220042204200422041;
defparam prom_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000002;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[29:0],dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 2;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h3CF000F03CE000E03000D00F600C0D20C0FCEE0F0E30D0E0D3034309700C0003;
defparam prom_inst_2.INIT_RAM_01 = 256'h00000C00000C0000D000080000000081028000000000000203B0E837C8300300;
defparam prom_inst_2.INIT_RAM_02 = 256'h02000000C2AC00000000808000000008C00000000C040C000002641080C040C0;
defparam prom_inst_2.INIT_RAM_03 = 256'h0000000000000A0000080020A20004C0200003000C2230040090004C00000000;
defparam prom_inst_2.INIT_RAM_04 = 256'h00000D0C010E300E20C030030010040003C00C00C002F2B20000000000300000;
defparam prom_inst_2.INIT_RAM_05 = 256'h300C3300C3300C30000000020000000000300000008000002000100010000000;
defparam prom_inst_2.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000003;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h34E000D034E000D03000F00EE00D4C50D040F10C0430C0C043030129332C0001;
defparam prom_inst_3.INIT_RAM_01 = 256'h00000C00000C0000F0000C00000000C303C000000000000243C0E03ECC300300;
defparam prom_inst_3.INIT_RAM_02 = 256'h02000000C154000000008000000000554000000000000C0000001020C00000C0;
defparam prom_inst_3.INIT_RAM_03 = 256'h0000000000000F00400C0030F30008803030C0000C2210080080000C20020000;
defparam prom_inst_3.INIT_RAM_04 = 256'h00000E0C020D310D30C030034010040000000C00C003C3C30000000000300000;
defparam prom_inst_3.INIT_RAM_05 = 256'h300C3300C3300C33000000030000000000200000008000002000200020002000;
defparam prom_inst_3.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000003;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[29:0],dout[9:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 2;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'h202820080028200808803A82EA0002200080320008082000808002840A2A0082;
defparam prom_inst_4.INIT_RAM_01 = 256'h2A08AA888200082200802A22222202880A008220822AAAA8EA754EAF1E228028;
defparam prom_inst_4.INIT_RAM_02 = 256'hA98AA08AA9588888888A8A8A08A08AD588888888A8A8AC22822B54128A8A8AC2;
defparam prom_inst_4.INIT_RAM_03 = 256'h22A2AAA22082252282260890E108AAAAA2A24A2A02919A26886222AA9A218888;
defparam prom_inst_4.INIT_RAM_04 = 256'hAAAA82000A020202102A0080A8AA2A2AAA88AC22480A23A108888208AA9A2A22;
defparam prom_inst_4.INIT_RAM_05 = 256'h020000200002000AA2A2080A08A08AAA28A08AA8A2822AAAA08AA08AA08AA08A;
defparam prom_inst_4.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000080;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[29:0],dout[11:10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 2;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h3104880E0105880604D816104580112808C112808C451808C42023000034304F;
defparam prom_inst_5.INIT_RAM_01 = 256'h84821E12038222080620318488488320E002208A20855560C9100C9100702086;
defparam prom_inst_5.INIT_RAM_02 = 256'h14E15821E002222222212121821821C0222222221212120860870048E1212120;
defparam prom_inst_5.INIT_RAM_03 = 256'h88385584822080486083820F08821DD838382087820C448123384825448CE122;
defparam prom_inst_5.INIT_RAM_04 = 256'h5556108123804480881842201202838560121A08220C0C088212088216048484;
defparam prom_inst_5.INIT_RAM_05 = 256'h468204782046820048486220A2122158820E21620818858446204E2046204E21;
defparam prom_inst_5.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000020;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[29:0],dout[13:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 2;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'h308444A9208444AD2044A448844809B4A4C09B4A4C2484A4C212934004B51243;
defparam prom_inst_6.INIT_RAM_01 = 256'h40410C41014911040110014044044012D09D104D10400004D59A8D59A9321241;
defparam prom_inst_6.INIT_RAM_02 = 256'h06904410C421111111101010410410C21111111101010104104309E490101010;
defparam prom_inst_6.INIT_RAM_03 = 256'h44A4101041104004104A41238E410CC1343410414846404011A4045440469011;
defparam prom_inst_6.INIT_RAM_04 = 256'h000048481348224AE481211201004A41040101041100AE2E4101044100404040;
defparam prom_inst_6.INIT_RAM_05 = 256'h254922549225492404041112910110014529100514B440156D1169116D116910;
defparam prom_inst_6.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000052;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[29:0],dout[15:14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 2;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'h79F455E179F455E17405F55FF45E9D85E5E9D85E5E75C5E5E717977FF7F59E77;
defparam prom_inst_7.INIT_RAM_01 = 256'h54515D51405D5545A5540D54554550D61781545154555557C1DFFC1DFD701755;
defparam prom_inst_7.INIT_RAM_02 = 256'h56155515D6ED555555551515515515EED5555555515151455457B83515151514;
defparam prom_inst_7.INIT_RAM_03 = 256'h5585555451545A4514585160F3515DD5F5F5D7545D6664591585450564561515;
defparam prom_inst_7.INIT_RAM_04 = 256'h55555C5D175E735E35D571579170585556914145D543E3E35151455155645454;
defparam prom_inst_7.INIT_RAM_05 = 256'h705D7705D7705D76454555561551555555615555558555556155615561556155;
defparam prom_inst_7.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000057;

endmodule //Gowin_pROM
